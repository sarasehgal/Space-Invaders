module InstantiateInvaders(
    input  logic        reset_ah, 
    input  logic        vsync,
    input  logic [7:0]  keycode,
    input  logic [9:0]  ShotX,
    input  logic [9:0]  ShotY,
    input  logic [9:0]  ShotW,
    input  logic [9:0]  ShotH,
    input  logic [49:0] Collision,

    output logic [9:0]  InvaderX[50], 
    output logic [9:0]  InvaderY[50],
    output logic [49:0] InvaderOn
    );
    logic col[10];
    logic [5:0] First_Active_Col;
    logic [5:0] Last_Active_Col;
    logic [3:0] Delay;
    
    always_comb begin
        col[0] = InvaderOn[0] | InvaderOn[10] | InvaderOn[20] | InvaderOn[30] | InvaderOn[40];
        col[1] = InvaderOn[1] | InvaderOn[11] | InvaderOn[21] | InvaderOn[31] | InvaderOn[41];
        col[2] = InvaderOn[2] | InvaderOn[12] | InvaderOn[22] | InvaderOn[32] | InvaderOn[42];
        col[3] = InvaderOn[3] | InvaderOn[13] | InvaderOn[23] | InvaderOn[33] | InvaderOn[43];
        col[4] = InvaderOn[4] | InvaderOn[14] | InvaderOn[24] | InvaderOn[34] | InvaderOn[44];
        col[5] = InvaderOn[5] | InvaderOn[15] | InvaderOn[25] | InvaderOn[35] | InvaderOn[45];
        col[6] = InvaderOn[6] | InvaderOn[16] | InvaderOn[26] | InvaderOn[36] | InvaderOn[46];
        col[7] = InvaderOn[7] | InvaderOn[17] | InvaderOn[27] | InvaderOn[37] | InvaderOn[47];
        col[8] = InvaderOn[8] | InvaderOn[18] | InvaderOn[28] | InvaderOn[38] | InvaderOn[48];
        col[9] = InvaderOn[9] | InvaderOn[19] | InvaderOn[29] | InvaderOn[39] | InvaderOn[49];
        for(int i = 0; i < 10; i++) begin
            if (col[i]) begin
                First_Active_Col = i;
                break;
            end
        end

        for(int i = 9; i >= 0; i--) begin
            if (col[i]) begin
                Last_Active_Col = i;
                break;
            end
        end
    end
    
    InvaderSpeed Speed (
        .InvaderOn(InvaderOn),
        .Delay(Delay)
    );
    
    invader invader0(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(150),
        .Invader_Y_Start(120),
        .InvaderS(8),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(0),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[0]),
        .Delay(Delay),
        .InvaderX(InvaderX[0]),
        .InvaderY(InvaderY[0]),
        .InvaderOn(InvaderOn[0])
      );
     
     invader invader1(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(175),
        .Invader_Y_Start(120),
        .InvaderS(8),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(0),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[1]),
        .Delay(Delay),
        .InvaderX(InvaderX[1]), 
        .InvaderY(InvaderY[1]),
        .InvaderOn(InvaderOn[1])
     );
     
     invader invader2(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(200),
        .Invader_Y_Start(120),
        .InvaderS(8),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(0),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[2]),
        .Delay(Delay),
        .InvaderX(InvaderX[2]), 
        .InvaderY(InvaderY[2]),
        .InvaderOn(InvaderOn[2])
     );
     
     invader invader3(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(225),
        .Invader_Y_Start(120),
        .InvaderS(8),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(0),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[3]),
        .Delay(Delay),
        .InvaderX(InvaderX[3]), 
        .InvaderY(InvaderY[3]),
        .InvaderOn(InvaderOn[3])
     );
     
     invader invader4(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(250),
        .Invader_Y_Start(120),
        .InvaderS(8),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(0),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[4]),
        .Delay(Delay),
        .InvaderX(InvaderX[4]), 
        .InvaderY(InvaderY[4]),
        .InvaderOn(InvaderOn[4])
     );
     
     invader invader5(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(275),
        .Invader_Y_Start(120),
        .InvaderS(8),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(0),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[5]),
        .Delay(Delay),
        .InvaderX(InvaderX[5]), 
        .InvaderY(InvaderY[5]),
        .InvaderOn(InvaderOn[5])
     );
     
     invader invader6(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(300),
        .Invader_Y_Start(120),
        .InvaderS(8),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(0),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[6]),
        .Delay(Delay),
        .InvaderX(InvaderX[6]), 
        .InvaderY(InvaderY[6]),
        .InvaderOn(InvaderOn[6])
     );
     
     invader invader7(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(325),
        .Invader_Y_Start(120),
        .InvaderS(8),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(0),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[7]),
        .Delay(Delay),
        .InvaderX(InvaderX[7]), 
        .InvaderY(InvaderY[7]),
        .InvaderOn(InvaderOn[7])
     );
     
     invader invader8(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(350),
        .Invader_Y_Start(120),
        .InvaderS(8),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(0),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[8]),
        .Delay(Delay),
        .InvaderX(InvaderX[8]), 
        .InvaderY(InvaderY[8]),
        .InvaderOn(InvaderOn[8])
     );
     
     invader invader9(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(375),
        .Invader_Y_Start(120),
        .InvaderS(8),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(0),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[9]),
        .Delay(Delay),
        .InvaderX(InvaderX[9]), 
        .InvaderY(InvaderY[9]),
        .InvaderOn(InvaderOn[9])
     );
     
    invader invader10(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(150),
        .Invader_Y_Start(145),
        .InvaderS(9),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(1),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[10]),
        .Delay(Delay),
        .InvaderX(InvaderX[10]),
        .InvaderY(InvaderY[10]),
        .InvaderOn(InvaderOn[10])
      );
     
     invader invader11(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(175),
        .Invader_Y_Start(145),
        .InvaderS(9),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(1),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[11]),
        .Delay(Delay),
        .InvaderX(InvaderX[11]), 
        .InvaderY(InvaderY[11]),
        .InvaderOn(InvaderOn[11])
     );
     
     invader invader12(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(200),
        .Invader_Y_Start(145),
        .InvaderS(9),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(1),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[12]),
        .Delay(Delay),
        .InvaderX(InvaderX[12]), 
        .InvaderY(InvaderY[12]),
        .InvaderOn(InvaderOn[12])
     );
     
     invader invader13(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(225),
        .Invader_Y_Start(145),
        .InvaderS(9),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(1),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[13]),
        .Delay(Delay),
        .InvaderX(InvaderX[13]), 
        .InvaderY(InvaderY[13]),
        .InvaderOn(InvaderOn[13])
     );
     
     invader invader14(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(250),
        .Invader_Y_Start(145),
        .InvaderS(9),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(1),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[14]),
        .Delay(Delay),
        .InvaderX(InvaderX[14]), 
        .InvaderY(InvaderY[14]),
        .InvaderOn(InvaderOn[14])
     );
     
     invader invader15(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(275),
        .Invader_Y_Start(145),
        .InvaderS(9),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(1),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[15]),
        .Delay(Delay),
        .InvaderX(InvaderX[15]), 
        .InvaderY(InvaderY[15]),
        .InvaderOn(InvaderOn[15])
     );
     
     invader invader16(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(300),
        .Invader_Y_Start(145),
        .InvaderS(9),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(1),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[16]),
        .Delay(Delay),
        .InvaderX(InvaderX[16]), 
        .InvaderY(InvaderY[16]),
        .InvaderOn(InvaderOn[16])
     );
     
     invader invader17(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(325),
        .Invader_Y_Start(145),
        .InvaderS(9),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(1),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[17]),
        .Delay(Delay),
        .InvaderX(InvaderX[17]), 
        .InvaderY(InvaderY[17]),
        .InvaderOn(InvaderOn[17])
     );
     
     invader invader18(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(350),
        .Invader_Y_Start(145),
        .InvaderS(9),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(1),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[18]),
        .Delay(Delay),
        .InvaderX(InvaderX[18]), 
        .InvaderY(InvaderY[18]),
        .InvaderOn(InvaderOn[18])
     );
     
     invader invader19(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(375),
        .Invader_Y_Start(145),
        .InvaderS(9),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(1),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[19]),
        .Delay(Delay),
        .InvaderX(InvaderX[19]), 
        .InvaderY(InvaderY[19]),
        .InvaderOn(InvaderOn[19])
     );
     
         invader invader20(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(150),
        .Invader_Y_Start(170),
        .InvaderS(9),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(2),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[20]),
        .Delay(Delay),
        .InvaderX(InvaderX[20]),
        .InvaderY(InvaderY[20]),
        .InvaderOn(InvaderOn[20])
      );
     
     invader invader21(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(175),
        .Invader_Y_Start(170),
        .InvaderS(9),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(2),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[21]),
        .Delay(Delay),
        .InvaderX(InvaderX[21]), 
        .InvaderY(InvaderY[21]),
        .InvaderOn(InvaderOn[21])
     );
     
     invader invader22(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(200),
        .Invader_Y_Start(170),
        .InvaderS(9),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(2),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[22]),
        .Delay(Delay),
        .InvaderX(InvaderX[22]), 
        .InvaderY(InvaderY[22]),
        .InvaderOn(InvaderOn[22])
     );
     
     invader invader23(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(225),
        .Invader_Y_Start(170),
        .InvaderS(9),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(2),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[23]),
        .Delay(Delay),
        .InvaderX(InvaderX[23]), 
        .InvaderY(InvaderY[23]),
        .InvaderOn(InvaderOn[23])
     );
     
     invader invader24(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(250),
        .Invader_Y_Start(170),
        .InvaderS(9),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(2),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[24]),
        .Delay(Delay),
        .InvaderX(InvaderX[24]), 
        .InvaderY(InvaderY[24]),
        .InvaderOn(InvaderOn[24])
     );
     
     invader invader25(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(275),
        .Invader_Y_Start(170),
        .InvaderS(9),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(2),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[25]),
        .Delay(Delay),
        .InvaderX(InvaderX[25]), 
        .InvaderY(InvaderY[25]),
        .InvaderOn(InvaderOn[25])
     );
     
     invader invader26(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(300),
        .Invader_Y_Start(170),
        .InvaderS(9),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(2),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[26]),
        .Delay(Delay),
        .InvaderX(InvaderX[26]), 
        .InvaderY(InvaderY[26]),
        .InvaderOn(InvaderOn[26])
     );
     
     invader invader27(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(325),
        .Invader_Y_Start(170),
        .InvaderS(9),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(2),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[27]),
        .Delay(Delay),
        .InvaderX(InvaderX[27]), 
        .InvaderY(InvaderY[27]),
        .InvaderOn(InvaderOn[27])
     );
     
     invader invader28(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(350),
        .Invader_Y_Start(170),
        .InvaderS(9),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(2),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[28]),
        .Delay(Delay),
        .InvaderX(InvaderX[28]), 
        .InvaderY(InvaderY[28]),
        .InvaderOn(InvaderOn[28])
     );
     
     invader invader29(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(375),
        .Invader_Y_Start(170),
        .InvaderS(9),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(2),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[29]),
        .Delay(Delay),
        .InvaderX(InvaderX[29]), 
        .InvaderY(InvaderY[29]),
        .InvaderOn(InvaderOn[29])
     );
     
         invader invader30(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(150),
        .Invader_Y_Start(195),
        .InvaderS(10),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(3),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[30]),
        .Delay(Delay),
        .InvaderX(InvaderX[30]),
        .InvaderY(InvaderY[30]),
        .InvaderOn(InvaderOn[30])
      );
     
     invader invader31(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(175),
        .Invader_Y_Start(195),
        .InvaderS(10),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(3),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[31]),
        .Delay(Delay),
        .InvaderX(InvaderX[31]), 
        .InvaderY(InvaderY[31]),
        .InvaderOn(InvaderOn[31])
     );
     
     invader invader32(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(200),
        .Invader_Y_Start(195),
        .InvaderS(10),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(3),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[32]),
        .Delay(Delay),
        .InvaderX(InvaderX[32]), 
        .InvaderY(InvaderY[32]),
        .InvaderOn(InvaderOn[32])
     );
     
     invader invader33(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(225),
        .Invader_Y_Start(195),
        .InvaderS(10),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(3),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[33]),
        .Delay(Delay),
        .InvaderX(InvaderX[33]), 
        .InvaderY(InvaderY[33]),
        .InvaderOn(InvaderOn[33])
     );
     
     invader invader34(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(250),
        .Invader_Y_Start(195),
        .InvaderS(10),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(3),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[34]),
        .Delay(Delay),
        .InvaderX(InvaderX[34]), 
        .InvaderY(InvaderY[34]),
        .InvaderOn(InvaderOn[34])
     );
     
     invader invader35(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(275),
        .Invader_Y_Start(195),
        .InvaderS(10),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(3),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[35]),
        .Delay(Delay),
        .InvaderX(InvaderX[35]), 
        .InvaderY(InvaderY[35]),
        .InvaderOn(InvaderOn[35])
     );
     
     invader invader36(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(300),
        .Invader_Y_Start(195),
        .InvaderS(10),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(3),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[36]),
        .Delay(Delay),
        .InvaderX(InvaderX[36]), 
        .InvaderY(InvaderY[36]),
        .InvaderOn(InvaderOn[36])
     );
     
     invader invader37(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(325),
        .Invader_Y_Start(195),
        .InvaderS(10),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(3),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[37]),
        .Delay(Delay),
        .InvaderX(InvaderX[37]), 
        .InvaderY(InvaderY[37]),
        .InvaderOn(InvaderOn[37])
     );
     
     invader invader38(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(350),
        .Invader_Y_Start(195),
        .InvaderS(10),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(3),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[38]),
        .Delay(Delay),
        .InvaderX(InvaderX[38]), 
        .InvaderY(InvaderY[38]),
        .InvaderOn(InvaderOn[38])
     );
     
     invader invader39(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(375),
        .Invader_Y_Start(195),
        .InvaderS(10),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(3),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[39]),
        .Delay(Delay),
        .InvaderX(InvaderX[39]), 
        .InvaderY(InvaderY[39]),
        .InvaderOn(InvaderOn[39])
     );
     
         invader invader40(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(150),
        .Invader_Y_Start(220),
        .InvaderS(10),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(4),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[40]),
        .Delay(Delay),
        .InvaderX(InvaderX[40]),
        .InvaderY(InvaderY[40]),
        .InvaderOn(InvaderOn[40])
      );
     
     invader invader41(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(175),
        .Invader_Y_Start(220),
        .InvaderS(10),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(4),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[41]),
        .Delay(Delay),
        .InvaderX(InvaderX[41]), 
        .InvaderY(InvaderY[41]),
        .InvaderOn(InvaderOn[41])
     );
     
     invader invader42(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(200),
        .Invader_Y_Start(220),
        .InvaderS(10),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(4),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[42]),
        .Delay(Delay),
        .InvaderX(InvaderX[42]), 
        .InvaderY(InvaderY[42]),
        .InvaderOn(InvaderOn[42])
     );
     
     invader invader43(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(225),
        .Invader_Y_Start(220),
        .InvaderS(10),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(4),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[43]),
        .Delay(Delay),
        .InvaderX(InvaderX[43]), 
        .InvaderY(InvaderY[43]),
        .InvaderOn(InvaderOn[43])
     );
     
     invader invader44(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(250),
        .Invader_Y_Start(220),
        .InvaderS(10),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(4),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[44]),
        .Delay(Delay),
        .InvaderX(InvaderX[44]), 
        .InvaderY(InvaderY[44]),
        .InvaderOn(InvaderOn[44])
     );
     
     invader invader45(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(275),
        .Invader_Y_Start(220),
        .InvaderS(10),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(4),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[45]),
        .Delay(Delay),
        .InvaderX(InvaderX[45]), 
        .InvaderY(InvaderY[45]),
        .InvaderOn(InvaderOn[45])
     );
     
     invader invader46(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(300),
        .Invader_Y_Start(220),
        .InvaderS(10),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(4),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[46]),
        .Delay(Delay),
        .InvaderX(InvaderX[46]), 
        .InvaderY(InvaderY[46]),
        .InvaderOn(InvaderOn[46])
     );
     
     invader invader47(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(325),
        .Invader_Y_Start(220),
        .InvaderS(10),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(4),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[47]),
        .Delay(Delay),
        .InvaderX(InvaderX[47]), 
        .InvaderY(InvaderY[47]),
        .InvaderOn(InvaderOn[47])
     );
     
     invader invader48(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(350),
        .Invader_Y_Start(220),
        .InvaderS(10),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(4),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[48]),
        .Delay(Delay),
        .InvaderX(InvaderX[48]), 
        .InvaderY(InvaderY[48]),
        .InvaderOn(InvaderOn[48])
     );
     
     invader invader49(
        .Reset(reset_ah), 
        .frame_clk(vsync),
        .Invader_X_Start(375),
        .Invader_Y_Start(220),
        .InvaderS(10),
        .keycode(keycode),
        .ShotX(ShotX),
        .ShotY(ShotY),
        .ShotW(ShotW), 
        .ShotH(ShotH),
        .index(4),
        .First_Active_Col(First_Active_Col),
        .Last_Active_Col(Last_Active_Col),
        .Collision(Collision[49]),
        .Delay(Delay),
        .InvaderX(InvaderX[49]), 
        .InvaderY(InvaderY[49]),
        .InvaderOn(InvaderOn[49])
     );
     
endmodule
